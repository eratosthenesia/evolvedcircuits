* simulation de RC2
.control
tran 10n 10000n
write
.endc

* Spice netlister for gnetlist
R5 n4 n5 1k
V1 n0 0 dc 1 ac 2 pulse 0 1 10n 10n 100n 1u 2u
R4 n3 n4 1k
R3 n2 n3 5k
C5 n5 0 1n
R2 n1 n2 1K
C4 n4 0 1n
R1 n0 n1 1k
C3 n3 0 1n
C2 n2 0 1n
C1 n1 0 1n
I1 n5 0 DC 0.01mA
R6 0 n5 10k
.END
